library ieee;
use ieee.std_logic_1164.all;

entity latchRS is
    port(reset, set       :    in std_logic;
         q, q_bar         :    inout std_logic);
end latchRS;

architecture funcionality of latchRS is
begin
	q     <= reset nor q_bar;
	q_bar <= set nor q;
end funcionality;