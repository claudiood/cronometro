library ieee;
use ieee.std_logic_1164.all;

entity decoder is
    port(D, C, B, A         : in std_logic;
         a, b, c, d, e, f   : out std_logic);
end decoder;

architecture funcionality of decoder is
begin

end funcionality;

